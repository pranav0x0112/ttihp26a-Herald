VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO PRAWNS_ART
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 33.0 BY 8.3 ;
  SYMMETRY X Y ;

  OBS
    LAYER Metal5 ;
      RECT 0 0 33.0 8.3 ;
  END

END PRAWNS_ART

END LIBRARY
