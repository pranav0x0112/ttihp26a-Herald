VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO PRAWNS_ART
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 33.0 BY 8.3 ;
  SYMMETRY X Y ;

END PRAWNS_ART

END LIBRARY
