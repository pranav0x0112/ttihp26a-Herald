// Blackbox wrapper for prawns_art GDS macro
(* blackbox *)
module PRAWNS_ART (
  input wire clk,
  output wire alive
);
  // This is a hard macro - no RTL implementation
endmodule
