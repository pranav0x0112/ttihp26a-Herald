(* blackbox *) (* keep *)
module PRAWNS_ART ();
endmodule
