// Pure decorative GDS art macro - blackbox only

`default_nettype none

(* blackbox *)
module PRAWNS_ART ();
endmodule
